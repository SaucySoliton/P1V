// top

/*
-------------------------------------------------------------------------------

This file is part of the hardware description for the Propeller 1 Design.

The Propeller 1 Design is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by the
Free Software Foundation, either version 3 of the License, or (at your option)
any later version.

The Propeller 1 Design is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
more details.

You should have received a copy of the GNU General Public License along with
the Propeller 1 Design.  If not, see <http://www.gnu.org/licenses/>.
-------------------------------------------------------------------------------
*/


`include "tim.v"
`include "dig.v"

module              top_veri
(
input               clock,           // clock input
input               inp_resn,           // reset input (active low)

inout       [31:0]  io,                 // i/o pins
input               sda_in,

output       [7:0]  ledg                // cog leds
);

`include "features.v"

//
// reg and wire declarations
//
reg                 nres;
wire         [7:0]  cfg;
wire        [31:0]  pin_out, pin_dir;
//wire                clkfb, clock_160, clk;
reg         [23:0]  reset_cnt;
reg                 reset_to;
wire                clk_pll;
wire                clk_cog;

wire         [31:0] pin_in = io;
assign              pin_in[28:0]=io[28:0];
assign              pin_in[31:30]=io[31:30];
assign              pin_in[29]=io[29]&sda_in;// Just a hack until we find the right way to do pullps
//    
// Clock control
//

tim clkgen( .clk        (clock),
            .res        (~inp_resn),
            .cfg        (cfg[6:0]),
            .clk_pll    (clk_pll),
            .clk_cog    (clk_cog)
          );

//
// Propeller 1 core module
//

dig core (  .nres       (nres),
            .cfg        (cfg),
            .clk_cog    (clk_cog),
            .clk_pll    (clk_pll),
            .pin_in     (pin_in),
            .pin_out    (pin_out),
            .pin_dir    (pin_dir),
            .cog_led    (ledg) );

always @ (posedge clk_cog)
    nres <= inp_resn & !cfg[7];

//
// Bidir I/O buffers
//

genvar i;
generate
    for (i=0; i<28; i=i+1)
    begin : iogen
        assign io[i] = pin_dir[i] ? pin_out[i] : 1'bZ;
    end
endgenerate

        assign io[28] = pin_dir[28] ? pin_out[28] : 1'b1;// I2C pullups
        assign io[29] = pin_dir[29] ? pin_out[29] : 1'b1;

        assign io[30] = pin_dir[30] ? pin_out[30] : 1'bZ;// Finish the rest
        assign io[31] = pin_dir[31] ? pin_out[31] : 1'bZ;


endmodule
